`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 08.10.2018 07:08:21
// Design Name: 
// Module Name: Control
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

/*
module Control(PNDNG, Ejecute,Lectura_Escritura,Hit,Desalojo,CLK,
                 Clear_Main_REG,Eneable_Main_REG, Sel_Mux_Bank,Eneable_REG, Clear_LDG_REG, Write_Eneable,
                 Banks_Eneable,R_W, Clear_Formador, Eneable_Formador,Sel_Mem_Mux);
input PNDNG, Ejecute,Lectura_Escritura,Hit,Desalojo, CLK;
output  Clear_Main_REG,Eneable_Main_REG, Sel_Mux_Bank,Eneable_REG;
output Clear_LDG_REG, Write_Eneable, Banks_Eneable,R_W, Clear_Formador, Eneable_Formador;
output [1:0]Sel_Mem_Mux;

Reg [12:0]OC  //Outputs Control

//always @(posedge CLK) begin

    //case({PNDNG, Ejecute,Lectura_Escritura,Hit,Desalojo,OC})
    
      //  default:
        
    
    
    //endcase

//end



endmodule

*/